//------------------------------------------------------------------------------
    //
    //  Filename       : fft_core.v
    //  Author         : liuxun
    //  Created        : 2019-12-03
    //  Description    : Fetch Wn for FFT
    //
//------------------------------------------------------------------------------

module fft_fetch_wn();

//*** PARAMETER ****************************************************************


//*** INPUT/OUTPUT *************************************************************


//*** WIRE/REG *****************************************************************


//*** MAIN BODY ****************************************************************



endmodule
