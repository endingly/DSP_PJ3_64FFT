//------------------------------------------------------------------------------
    //
    //  Filename       : fft_fetch_data.v
    //  Author         : liuxun
    //  Created        : 2019-12-03
    //  Description    : Fetch 64 re and im data for FFT
    //                   and do reorder as well.
//------------------------------------------------------------------------------

`include "../include/fft_defines.vh"

module fft_fetch_data();

//*** PARAMETER ****************************************************************


//*** INPUT/OUTPUT *************************************************************


//*** WIRE/REG *****************************************************************


//*** MAIN BODY ****************************************************************


endmodule
