//------------------------------------------------------------------------------
    //
    //  Filename       : fft_top.v
    //  Author         : liuxun
    //  Created        : 2019-12-03
    //  Description    : Build FFT using fft_core2 module with a pipeline of 6
    //
//------------------------------------------------------------------------------

`include "../include/fft_defines.vh"
module fft_top();

//*** PARAMETER ****************************************************************


//*** INPUT/OUTPUT *************************************************************


//*** WIRE/REG *****************************************************************


//*** MAIN BODY ****************************************************************



endmodule
